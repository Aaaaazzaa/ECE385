//module audio_toplevel(
//  input logic CLOCK_50,
//  input	logic	CLOCK_27,
//	// Avalon Reset Input
//	input logic RESET,
//  input	logic	[3:0]	KEY,
//  input	logic	[3:0]	SW,
//  input	logic			AUD_ADCDAT,
//  // Bidirectionals
//  inout	logic 			AUD_BCLK,
//  inout	logic			AUD_ADCLRCK,
//  inout	logic	AUD_DACLRCK,
//  inout	logic	I2C_SDAT,
//  // Outputs
//  output logic	AUD_XCK,
//  output logic	AUD_DACDAT,
//  output logic	I2C_SCLK,
//  output 		[6:0] HEX0, HEX1, HEX2, HEX3, HEX4, HEX4, HEX5, HEX6, HEX7,
//  output 		[8:0] LEDG,
//  output logic [12:0] DRAM_ADDR,
//  output logic [1:0]  DRAM_BA,
//  output logic        DRAM_CAS_N,
//  output logic        DRAM_CKE,
//  output logic        DRAM_CS_N,
//  inout  logic [31:0] DRAM_DQ,
//  output logic [3:0]  DRAM_DQM,
//  output logic        DRAM_RAS_N,
//  output logic        DRAM_WE_N,
//  output logic        DRAM_CLK
//  );
//
//
//
//
//endmodule
