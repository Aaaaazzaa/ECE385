module test(input logic [9:0] register [3],
				output logic [1:0] whatever);
assign whatever = 2'd10/2'd2;
endmodule 