module audio_controller