// Copyright (C) 2018  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details.

// Generated by Quartus Prime Version 18.0.0 Build 614 04/24/2018 SJ Lite Edition
// Created on Sat Feb 09 15:28:22 2019

// synthesis message_off 10175

`timescale 1ns/1ns

module state_machine (
    input reset, input clock, input Reset, input Exe,
    output Add);

    enum int unsigned { S1=0, S2=1, S0=2, start_reset=3, S3=4, S4=5, S5=6, S6=7, S7Add=8, halt=9 } fstate, reg_fstate;

    always_ff @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always_comb begin
        if (reset) begin
            reg_fstate <= start_reset;
            Add <= 1'b0;
        end
        else begin
            Add <= 1'b0;
            case (fstate)
                S1: begin
                    if (~(Reset))
                        reg_fstate <= S2;
                    else if (Reset)
                        reg_fstate <= start_reset;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= S1;

                    if ((Exe == 1'b1))
                        Add <= 1'b1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        Add <= 1'b0;
                end
                S2: begin
                    if (~(Reset))
                        reg_fstate <= S3;
                    else if (Reset)
                        reg_fstate <= start_reset;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= S2;
                end
                S0: begin
                    if (~(Reset))
                        reg_fstate <= S1;
                    else if (Reset)
                        reg_fstate <= start_reset;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= S0;
                end
                start_reset: begin
                    if ((~(Reset) & Exe))
                        reg_fstate <= S0;
                    else if (((Reset & Exe) | ~(Exe)))
                        reg_fstate <= start_reset;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= start_reset;
                end
                S3: begin
                    if (~(Reset))
                        reg_fstate <= S4;
                    else if (Reset)
                        reg_fstate <= start_reset;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= S3;
                end
                S4: begin
                    if (~(Reset))
                        reg_fstate <= S5;
                    else if (Reset)
                        reg_fstate <= start_reset;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= S4;
                end
                S5: begin
                    if (~(Reset))
                        reg_fstate <= S6;
                    else if (Reset)
                        reg_fstate <= halt;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= S5;
                end
                S6: begin
                    if (~(Reset))
                        reg_fstate <= S7Add;
                    else if (Reset)
                        reg_fstate <= start_reset;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= S6;
                end
                S7Add: begin
                    if (~(Reset))
                        reg_fstate <= halt;
                    else if (Reset)
                        reg_fstate <= start_reset;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= S7Add;
                end
                halt: begin
                    if ((Reset | ~(Exe)))
                        reg_fstate <= start_reset;
                    else if ((Exe & ~(Reset)))
                        reg_fstate <= halt;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= halt;
                end
                default: begin
                    Add <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // state_machine
