module stateISB(  input state,
                  output result);





endmodule
