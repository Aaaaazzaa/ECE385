// Copyright (C) 2018  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details.

// Generated by Quartus Prime Version 18.0.0 Build 614 04/24/2018 SJ Lite Edition
// Created on Sat Apr 20 22:15:47 2019

// synthesis message_off 10175

`timescale 1ns/1ns

module adc_sm (
    input logic reset, input logic clock, input logic INIT_FINISH, input logic adc_full,
    output logic INIT);

    enum int unsigned { Init=0, Gather=1, Store=2 } fstate, reg_fstate;

    always_ff @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always_comb begin
        if (reset) begin
            reg_fstate <= Init;
            INIT <= 1'b0;
        end
        else begin
            INIT <= 1'b0;
            case (fstate)
                Init: begin
                    if (INIT_FINISH)
                        reg_fstate <= Gather;
                    else if (~(INIT_FINISH))
                        reg_fstate <= Init;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= Init;

                    INIT <= 1'b1;
                end
                Gather: begin
                    if (adc_full)
                        reg_fstate <= Store;
                    else if (~(adc_full))
                        reg_fstate <= Gather;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= Gather;
                end
                Store: begin
                    if (~(adc_full))
                        reg_fstate <= Gather;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= Store;
                end
                default: begin
                    INIT <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // adc_sm
