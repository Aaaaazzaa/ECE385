// Copyright (C) 2018  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details.

// Generated by Quartus Prime Version 18.0.0 Build 614 04/24/2018 SJ Lite Edition
// Created on Mon Apr 15 18:51:05 2019

// synthesis message_off 10175

`timescale 1ns/1ns

module sramcontroller (
    input reset, input clock, input ReadDone, input Blank,
    output Clear, output BufferWE, output UpdateAddr);

    enum int unsigned { ReadOnly=0, ClearFrame=1, SetAddr=2, WaitSRAM=3, EndOfNotch=4 } fstate, reg_fstate;

    always_ff @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always_comb begin
        if (reset) begin
            reg_fstate <= ClearFrame;
            Clear <= 1'b0;
            BufferWE <= 1'b0;
            UpdateAddr <= 1'b0;
        end
        else begin
            Clear <= 1'b0;
            BufferWE <= 1'b0;
            UpdateAddr <= 1'b0;
            case (fstate)
                ReadOnly: begin
                    if (~(Blank))
                        reg_fstate <= ClearFrame;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= ReadOnly;

                    BufferWE <= 1'b1;
                end
                ClearFrame: begin
                    reg_fstate <= SetAddr;

                    Clear <= 1'b1;
                end
                SetAddr: begin
                    reg_fstate <= WaitSRAM;
                end
                WaitSRAM: begin
                    if (~(ReadDone))
                        reg_fstate <= SetAddr;
                    else if (ReadDone)
                        reg_fstate <= EndOfNotch;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= WaitSRAM;

                    UpdateAddr <= 1'b1;
                end
                EndOfNotch: begin
                    if (Blank)
                        reg_fstate <= ReadOnly;
                    else if (~(Blank))
                        reg_fstate <= EndOfNotch;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= EndOfNotch;
                end
                default: begin
                    Clear <= 1'bx;
                    BufferWE <= 1'bx;
                    UpdateAddr <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // SM1
