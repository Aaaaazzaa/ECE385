    Mac OS X            	   2  �     �                                    ATTR;���  �  $  l                 $   9  com.apple.quarantine   ]     com.apple.lastuseddate#PS 36-  m   5  )com.apple.metadata:kMDItemDownloadedDate   �   �  %com.apple.metadata:kMDItemWhereFroms 0083;5c94344c;Safari;54F8644C-B66B-4B36-A100-48639D312BCB�4�\    �I>    bplist00�3A�"5�oU�
                            bplist00�_{https://wiki.illinois.edu/wiki/download/attachments/688237958/audio_interface.vhd?version=1&modificationDate=1547245710000&_?https://wiki.illinois.edu/wiki/display/ece385sp19/Final+Project�                            �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               This resource fork intentionally left blank                                                                                                                                                                                                                            ��