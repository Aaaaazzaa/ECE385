// Copyright (C) 2018  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details.

// Generated by Quartus Prime Version 18.0.0 Build 614 04/24/2018 SJ Lite Edition
// Created on Fri Feb 15 14:46:42 2019

// synthesis message_off 10175

`timescale 1ns/1ns

module state (
    input logic reset, input logic clock, input logic  M, input logic Exe,
    output logic Shift, output logic Add, output logic  Sub, output logic Clr_Ld);

    enum int unsigned { Start=0, S0=1, S1=2, S2=3, S3=4, S4=5, S5=6, S6=7, S7=8, Halt=9, Add0=10, Add1=11, Add2=12, Add3=13, Add4=14, Add5=15, Add6=16, Sub7=17, S8=18, Display=19 } fstate, reg_fstate;

    always_ff @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always_comb begin
        if (reset) begin
            reg_fstate <= Display;
            Shift <= 1'b0;
            Add <= 1'b0;
            Sub <= 1'b0;
            Clr_Ld <= 1'b0;
        end
        else begin
            Shift <= 1'b0;
            Add <= 1'b0;
            Sub <= 1'b0;
            Clr_Ld <= 1'b0;
            case (fstate)
                Start: begin
                    reg_fstate <= S0;

                    Clr_Ld <= 1'b1;
                end
                S0: begin
                    if (~(M))
                        reg_fstate <= S1;
                    else if (M)
                        reg_fstate <= Add0;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= S0;

                    Shift <= 1'b1;
                end
                S1: begin
                    if (~(M))
                        reg_fstate <= S2;
                    else if (M)
                        reg_fstate <= Add1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= S1;

                    Shift <= 1'b1;
                end
                S2: begin
                    if (~(M))
                        reg_fstate <= S3;
                    else if (M)
                        reg_fstate <= Add2;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= S2;

                    Shift <= 1'b1;
                end
                S3: begin
                    if (~(M))
                        reg_fstate <= S4;
                    else if (M)
                        reg_fstate <= Add3;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= S3;

                    Shift <= 1'b1;
                end
                S4: begin
                    if (~(M))
                        reg_fstate <= S5;
                    else if (M)
                        reg_fstate <= Add4;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= S4;

                    Shift <= 1'b1;
                end
                S5: begin
                    if (~(M))
                        reg_fstate <= S6;
                    else if (M)
                        reg_fstate <= Add5;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= S5;

                    Shift <= 1'b1;
                end
                S6: begin
                    if (~(M))
                        reg_fstate <= S7;
                    else if (M)
                        reg_fstate <= Add6;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= S6;

                    Shift <= 1'b1;
                end
                S7: begin
                    if (M)
                        reg_fstate <= Sub7;
                    else if (~(M))
                        reg_fstate <= S8;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= S7;

                    Shift <= 1'b1;
                end
                Halt: begin
                    if (~(Exe))
                        reg_fstate <= Display;
                    else if (Exe)
                        reg_fstate <= Halt;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= Halt;
                end
                Add0: begin
                    reg_fstate <= S1;

                    Add <= 1'b1;
                end
                Add1: begin
                    reg_fstate <= S2;

                    Add <= 1'b1;
                end
                Add2: begin
                    reg_fstate <= S3;

                    Add <= 1'b1;
                end
                Add3: begin
                    reg_fstate <= S4;

                    Add <= 1'b1;
                end
                Add4: begin
                    reg_fstate <= S5;

                    Add <= 1'b1;
                end
                Add5: begin
                    reg_fstate <= S6;

                    Add <= 1'b1;
                end
                Add6: begin
                    reg_fstate <= S7;

                    Add <= 1'b1;
                end
                Sub7: begin
                    reg_fstate <= S8;

                    Sub <= 1'b1;
                end
                S8: begin
                    reg_fstate <= Halt;

                    Shift <= 1'b1;
                end
                Display: begin
                    if (Exe)
                        reg_fstate <= Start;
                    else if (~(Exe))
                        reg_fstate <= Display;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= Display;
                end
                default: begin
                    Shift <= 1'bx;
                    Add <= 1'bx;
                    Sub <= 1'bx;
                    Clr_Ld <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // state
