module colorMapper();


endmodule 