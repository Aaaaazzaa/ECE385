module Control(	input logic Reset, Clk, Run, ClearA_LoadB,
						output logic Clr_Ld, Shift, Add, Sub);
						
						
						
						
						
						
						
						
						
						
						
						
						
						
						
endmodule 