//module unpacked(input Clk, Reset,
//							output A00);
//							
//		logic [3:0] A [50000];
//		always_ff @ (posedge Clk) begin
//			if (Reset)
//				A <= 20000'b0;
//			end
//		assign A00 = A[0][0];
//							
//							
//endmodule
							