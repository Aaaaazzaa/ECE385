// Copyright (C) 2018  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions
// and other software and tools, and its AMPP partner logic
// functions, and any output files from any of the foregoing
// (including device programming or simulation files), and any
// associated documentation or information are expressly subject
// to the terms and conditions of the Intel Program License
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details.

// Generated by Quartus Prime Version 18.0.0 Build 614 04/24/2018 SJ Lite Edition
// Created on Sun Apr 21 15:21:29 2019

// synthesis message_off 10175

`timescale 1ns/1ns

module convolutionSM (
    input  logic reset, input  logic clock, input  logic interDone, input  logic arrDone, input  logic inBlock,
    output  logic nUpdate, output logic  Clear, output  logic Done, output logic  mUpdate, output logic  store);

    enum int unsigned { interLoop=0, arrLoop=1, Start=2, Idle=3, singleStore=4 } fstate, reg_fstate;

    always_ff @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always_comb begin
        if (reset) begin
            reg_fstate <= Start;
            nUpdate <= 1'b0;
            Clear <= 1'b0;
            Done <= 1'b0;
            mUpdate <= 1'b0;
            store <= 1'b0;
        end
        else begin
            nUpdate <= 1'b0;
            Clear <= 1'b0;
            Done <= 1'b0;
            mUpdate <= 1'b0;
            store <= 1'b0;
            case (fstate)
                interLoop: begin
                    if (interDone)
                        reg_fstate <= singleStore;
                    else if (~(interDone))
                        reg_fstate <= interLoop;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= interLoop;

                    mUpdate <= 1'b1;
                end
                arrLoop: begin
                    if (~(arrDone))
                        reg_fstate <= interLoop;
                    else if (arrDone)
                        reg_fstate <= Idle;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= arrLoop;

                    Clear <= 1'b1;

                    nUpdate <= 1'b1;
                end
                Start: begin
                    reg_fstate <= arrLoop;
                end
                Idle: begin
                    if (~(inBlock))
                        reg_fstate <= Start;
                    else if (inBlock)
                        reg_fstate <= Idle;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= Idle;

                    Done <= 1'b1;
                end
                singleStore: begin
                    reg_fstate <= arrLoop;

                    store <= 1'b1;
                end
                default: begin
                    nUpdate <= 1'bx;
                    Clear <= 1'bx;
                    Done <= 1'bx;
                    mUpdate <= 1'bx;
                    store <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // convolutionSM
