module terrain( );




endmodule
