// Copyright (C) 2018  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details.

// Generated by Quartus Prime Version 18.0.0 Build 614 04/24/2018 SJ Lite Edition
// Created on Fri Apr 19 17:26:43 2019

// synthesis message_off 10175

`timescale 1ns/1ns

module convolution (
    input logic reset, input logic clock, input logic counter, input logic start,
    output logic Convolve);

    enum int unsigned { Finished=0, Start=1, Convolution=2 } fstate, reg_fstate;

    always_ff @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always_comb begin
        if (reset) begin
            reg_fstate <= Start;
            Convolve <= 1'b0;
        end
        else begin
            Convolve <= 1'b0;
            case (fstate)
                Finished: begin
                    reg_fstate <= Start;

                    Convolve <= 1'b0;
                end
                Start: begin
                    if (start)
                        reg_fstate <= Convolution;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= Start;

                    Convolve <= 1'b0;
                end
                Convolution: begin
                    if (~(counter))
                        reg_fstate <= Finished;
                    else if (counter)
                        reg_fstate <= Convolution;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= Convolution;

                    Convolve <= 1'b1;
                end
                default: begin
                    Convolve <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // convolution
