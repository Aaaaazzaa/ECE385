// Copyright (C) 2018  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions
// and other software and tools, and its AMPP partner logic
// functions, and any output files from any of the foregoing
// (including device programming or simulation files), and any
// associated documentation or information are expressly subject
// to the terms and conditions of the Intel Program License
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details.

// Generated by Quartus Prime Version 18.0.0 Build 614 04/24/2018 SJ Lite Edition
// Created on Fri Mar 29 20:32:22 2019

// synthesis message_off 10175

`timescale 1ns/1ns

module Lab9_mealy_sm (
    input logic reset, input logic clock, input logic AES_START, input logic Cycle, input logic IMCDone,
    output logic Update, output logic AES_DONE, output logic Clear, output logic SelL, output logic SelH, output logic Store, output logic UpdateIMC);

    enum int unsigned { ISB10=9, ARK10=10, Done=11, Reset=1, ISR10=8, Idle=0, ISR=3, ARK0=2, ISB=4, IMC=6, ARK=5, IMCWait=7 } fstate, reg_fstate;

    always_ff @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always_comb begin
        if (reset) begin
            reg_fstate <= Idle;
            Update <= 1'b0;
            AES_DONE <= 1'b0;
            Clear <= 1'b0;
            SelL <= 1'b0;
            SelH <= 1'b0;
            Store <= 1'b0;
            UpdateIMC <= 1'b0;
        end
        else begin
            Update <= 1'b0;
            AES_DONE <= 1'b0;
            Clear <= 1'b0;
            SelL <= 1'b0;
            SelH <= 1'b0;
            Store <= 1'b0;
            UpdateIMC <= 1'b0;
            case (fstate)
                ISB10: begin
                    reg_fstate <= ARK10;

                    SelL <= 1'b1;

                    Store <= 1'b1;
                end
                ARK10: begin
                    reg_fstate <= Done;

                    SelL <= 1'b0;

                    Store <= 1'b1;
                end
                Done: begin
                    if (~(AES_START))
                        reg_fstate <= Idle;
                    else if (AES_START)
                        reg_fstate <= Done;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= Done;

                    AES_DONE <= 1'b1;
                end
                Reset: begin
                    reg_fstate <= ARK0;

                    Clear <= 1'b1;
                end
                ISR10: begin
                    reg_fstate <= ISB10;

                    Store <= 1'b1;

                    SelH <= 1'b1;
                end
                Idle: begin
                    if (AES_START)
                        reg_fstate <= Reset;
                    else if (~(AES_START))
                        reg_fstate <= Idle;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= Idle;
                end
                ISR: begin
                    reg_fstate <= ISB;

                    Store <= 1'b1;

                    SelH <= 1'b1;
                end
                ARK0: begin
                    reg_fstate <= ISR;

                    SelL <= 1'b0;

                    Store <= 1'b1;

                    Update <= 1'b1;
                end
                ISB: begin
                    reg_fstate <= ARK;

                    SelL <= 1'b1;
                    SelL <= 1'b1;

                    Store <= 1'b1;
                end
                IMC: begin
                    if (IMCDone)
                        reg_fstate <= IMCWait;
                    else if (~(IMCDone))
                        reg_fstate <= IMC;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= IMC;

                    SelL <= 1'b0;

                    UpdateIMC <= 1'b1;

                    Store <= 1'b0;

                    SelH <= 1'b0;
                end
                ARK: begin
                    reg_fstate <= IMC;

                    SelL <= 1'b0;

                    Store <= 1'b1;

                    Update <= 1'b1;
                end
                IMCWait: begin
                    if (~(Cycle))
                        reg_fstate <= ISR10;
                    else if (Cycle)
                        reg_fstate <= ISR;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= IMCWait;

                    SelL <= 1'b1;

                    Store <= 1'b1;

                    SelH <= 1'b1;
                end
                default: begin
                    Update <= 1'bx;
                    AES_DONE <= 1'bx;
                    Clear <= 1'bx;
                    SelL <= 1'bx;
                    SelH <= 1'bx;
                    Store <= 1'bx;
                    UpdateIMC <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // Lab9_mealy_sm
